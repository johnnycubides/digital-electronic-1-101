module testbech;

  // STIMULUS
  // reg a = 0, b = 0;
  // initial
  // begin
  //   # 17 a = 1, b = 1;
  //   # 11 a = 1, b = 0;
  //   # 29 a = 1, b = 1;
  //   # 11 a = 1, b = 0;
  //   # 100 $finish(); // [stop(), $finish()]
  // end

  reg [2:0] inputs;
  // inputs[0] inputs[1] inputs[2]
  // integer i;
  // initial
  // begin
  //   for (i=0; i<8; i=i+1)
  //   begin
  //     inputs = i;
  //     #1;
  //   end
  // end

  // CLOCK STIMULUS
  // Make a regular pulsing clock.
  // reg clk = 0;
  // always #5 clk = !clk;

  // RESULT FOR DEVICE/DESIGN UNDER TEST
  wire [1:0] outs;
  // DEVICE/DESIGN UNDER TEST
  fulladder dut (
    .in_b(inputs[2]), .in_a(inputs[1]), .in_ci(inputs[0]),
    .out_co(outs[1]), .out_s(outs[0])
  );

  // STIMULUS ARGS
  initial
  begin
    if(! $value$plusargs("inputs=%b", inputs)) begin
      $display("ERROR: please specify +inputs=<value> to start.");
      $finish;
    end

    wait (outs) $display("outs = %d", outs);
    #1
    $finish;
  end

  // MONITOR
  // initial
  //   $monitor("Time: %t, a = %d, b = %d => out = %d",
  //     $time, a, b, value);

  // WAVES IN VCD TO OPEN IN GTKWAVE
  initial
  begin
    $dumpfile("top.vcd");
    $dumpvars(0, testbech);
  end


endmodule

module top(input b, a, cin, output cout, s);
fulladder fulladder(b,a,cin,cout,s);
endmodule

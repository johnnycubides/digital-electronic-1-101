module and3 (input a, b , c, output z);
  assign z = a & b & c;
endmodule

// 8N1 UART Module, transmit only

module uart_tx_8n1 (
    clk,  // input clock
    txbyte,  // outgoing byte
    senddata,  // trigger tx
    txdone,  // outgoing byte sent
    tx  // tx wire
);

  /* Inputs */
  input clk;
  input [7:0] txbyte;
  input senddata;

  /* Outputs */
  output txdone;
  output tx;

  /* Parameters */
  parameter STATE_IDLE = 8'd0;
  parameter STATE_STARTTX = 8'd1;
  parameter STATE_TXING = 8'd2;
  parameter STATE_TXDONE = 8'd3;

  /* State variables */
  reg [7:0] state = 8'b0;
  reg [7:0] buf_tx = 8'b0;
  reg [7:0] bits_sent = 8'b0;
  reg txbit = 1'b1;
  reg txdone = 1'b0;

  /* Wiring */
  assign tx = txbit;

  /* always */
  always @(posedge clk) begin
    // start sending?
    if (senddata == 1 && state == STATE_IDLE) begin
      state  <= STATE_STARTTX;
      buf_tx <= txbyte;
      txdone <= 1'b0;
    end else if (state == STATE_IDLE) begin
      // idle at high
      txbit  <= 1'b1;
      txdone <= 1'b0;
    end

    // send start bit (low)
    if (state == STATE_STARTTX) begin
      txbit <= 1'b0;
      state <= STATE_TXING;
    end
    // clock data out
    if (state == STATE_TXING && bits_sent < 8'd8) begin
      txbit  <= buf_tx[0];
      buf_tx <= buf_tx >> 1;
      bits_sent = bits_sent + 1;
    end else if (state == STATE_TXING) begin
      // send stop bit (high)
      txbit <= 1'b1;
      bits_sent <= 8'b0;
      state <= STATE_TXDONE;
    end

    // tx done
    if (state == STATE_TXDONE) begin
      txdone <= 1'b1;
      state  <= STATE_IDLE;
    end

  end

endmodule


module gate_or (input a, b, output c);
  assign c = a | b;
endmodule
